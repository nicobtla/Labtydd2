library verilog;
use verilog.vl_types.all;
entity partea_vlg_vec_tst is
end partea_vlg_vec_tst;
