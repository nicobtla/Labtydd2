library verilog;
use verilog.vl_types.all;
entity parteA_vlg_vec_tst is
end parteA_vlg_vec_tst;
