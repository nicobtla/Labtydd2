library verilog;
use verilog.vl_types.all;
entity parteb_vlg_vec_tst is
end parteb_vlg_vec_tst;
