library verilog;
use verilog.vl_types.all;
entity esquematico_vlg_check_tst is
    port(
        cout            : in     vl_logic;
        s1              : in     vl_logic;
        s2              : in     vl_logic;
        s3              : in     vl_logic;
        s4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end esquematico_vlg_check_tst;
