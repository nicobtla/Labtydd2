library verilog;
use verilog.vl_types.all;
entity SM1_vlg_vec_tst is
end SM1_vlg_vec_tst;
