library verilog;
use verilog.vl_types.all;
entity esquematico_vlg_vec_tst is
end esquematico_vlg_vec_tst;
