library verilog;
use verilog.vl_types.all;
entity sumador_completo_vlg_vec_tst is
end sumador_completo_vlg_vec_tst;
